library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;
--library unisim;
--use unisim.vcomponents.all;

entity square_drawer_tb is
  generic (
    -- Generics go here...
  );
  port (
    -- Inputs, outputs, inouts go here...
  );
end entity;


