-- soc_video_system.vhd

-- Generated using ACDS version 17.1 590

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity soc_video_system is
	port (
		clk_clk                          : in    std_logic                     := '0';             --              clk.clk
		clk_sdram_clk                    : out   std_logic;                                        --        clk_sdram.clk
		clk_video_clk                    : out   std_logic;                                        --        clk_video.clk
		edge_detect_bypass               : in    std_logic                     := '0';             --      edge_detect.bypass
		reset_reset_n                    : in    std_logic                     := '0';             --            reset.reset_n
		vga_CLK                          : out   std_logic;                                        --              vga.CLK
		vga_HS                           : out   std_logic;                                        --                 .HS
		vga_VS                           : out   std_logic;                                        --                 .VS
		vga_BLANK                        : out   std_logic;                                        --                 .BLANK
		vga_SYNC                         : out   std_logic;                                        --                 .SYNC
		vga_R                            : out   std_logic_vector(7 downto 0);                     --                 .R
		vga_G                            : out   std_logic_vector(7 downto 0);                     --                 .G
		vga_B                            : out   std_logic_vector(7 downto 0);                     --                 .B
		video_config_SDAT                : inout std_logic                     := '0';             --     video_config.SDAT
		video_config_SCLK                : out   std_logic;                                        --                 .SCLK
		video_in_decoder_PIXEL_CLK       : in    std_logic                     := '0';             -- video_in_decoder.PIXEL_CLK
		video_in_decoder_LINE_VALID      : in    std_logic                     := '0';             --                 .LINE_VALID
		video_in_decoder_FRAME_VALID     : in    std_logic                     := '0';             --                 .FRAME_VALID
		video_in_decoder_pixel_clk_reset : in    std_logic                     := '0';             --                 .pixel_clk_reset
		video_in_decoder_PIXEL_DATA      : in    std_logic_vector(11 downto 0) := (others => '0'); --                 .PIXEL_DATA
		video_merge_export               : in    std_logic                     := '0';             --      video_merge.export
		video_sdram_addr                 : out   std_logic_vector(12 downto 0);                    --      video_sdram.addr
		video_sdram_ba                   : out   std_logic_vector(1 downto 0);                     --                 .ba
		video_sdram_cas_n                : out   std_logic;                                        --                 .cas_n
		video_sdram_cke                  : out   std_logic;                                        --                 .cke
		video_sdram_cs_n                 : out   std_logic;                                        --                 .cs_n
		video_sdram_dq                   : inout std_logic_vector(15 downto 0) := (others => '0'); --                 .dq
		video_sdram_dqm                  : out   std_logic_vector(1 downto 0);                     --                 .dqm
		video_sdram_ras_n                : out   std_logic;                                        --                 .ras_n
		video_sdram_we_n                 : out   std_logic;                                        --                 .we_n
		video_split_export               : in    std_logic                     := '0'              --      video_split.export
	);
end entity soc_video_system;

architecture rtl of soc_video_system is
	component soc_video_system_altpll_0 is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component soc_video_system_altpll_0;

	component soc_video_system_audio_and_video_config_0 is
		port (
			clk         : in    std_logic                     := 'X';             -- clk
			reset       : in    std_logic                     := 'X';             -- reset
			address     : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			byteenable  : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			read        : in    std_logic                     := 'X';             -- read
			write       : in    std_logic                     := 'X';             -- write
			writedata   : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			readdata    : out   std_logic_vector(31 downto 0);                    -- readdata
			waitrequest : out   std_logic;                                        -- waitrequest
			I2C_SDAT    : inout std_logic                     := 'X';             -- export
			I2C_SCLK    : out   std_logic                                         -- export
		);
	end component soc_video_system_audio_and_video_config_0;

	component soc_video_system_fpga_only_master is
		generic (
			USE_PLI     : integer := 0;
			PLI_PORT    : integer := 50000;
			FIFO_DEPTHS : integer := 2
		);
		port (
			clk_clk              : in  std_logic                     := 'X';             -- clk
			clk_reset_reset      : in  std_logic                     := 'X';             -- reset
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_readdata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			master_read          : out std_logic;                                        -- read
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(31 downto 0);                    -- writedata
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_byteenable    : out std_logic_vector(3 downto 0);                     -- byteenable
			master_reset_reset   : out std_logic                                         -- reset
		);
	end component soc_video_system_fpga_only_master;

	component soc_video_system_pixel_buffer is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component soc_video_system_pixel_buffer;

	component soc_video_system_pixel_onchip_buffer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(17 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(7 downto 0);                     -- readdata
			writedata  : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component soc_video_system_pixel_onchip_buffer;

	component altera_up_avalon_video_edge_detection is
		generic (
			WIDTH : integer := 640
		);
		port (
			clk               : in  std_logic                    := 'X';             -- clk
			reset             : in  std_logic                    := 'X';             -- reset
			bypass            : in  std_logic                    := 'X';             -- bypass
			in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			in_valid          : in  std_logic                    := 'X';             -- valid
			in_ready          : out std_logic;                                       -- ready
			out_data          : out std_logic_vector(7 downto 0);                    -- data
			out_startofpacket : out std_logic;                                       -- startofpacket
			out_endofpacket   : out std_logic;                                       -- endofpacket
			out_valid         : out std_logic;                                       -- valid
			out_ready         : in  std_logic                    := 'X'              -- ready
		);
	end component altera_up_avalon_video_edge_detection;

	component soc_video_system_video_bayer_resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_data          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic                                         -- valid
		);
	end component soc_video_system_video_bayer_resampler;

	component soc_video_system_video_clipper is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_data          : out std_logic_vector(23 downto 0);                    -- data
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic                                         -- valid
		);
	end component soc_video_system_video_clipper;

	component soc_video_system_video_decoder_0 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                     -- data
			PIXEL_CLK                : in  std_logic                     := 'X';             -- export
			LINE_VALID               : in  std_logic                     := 'X';             -- export
			FRAME_VALID              : in  std_logic                     := 'X';             -- export
			pixel_clk_reset          : in  std_logic                     := 'X';             -- export
			PIXEL_DATA               : in  std_logic_vector(11 downto 0) := (others => 'X')  -- export
		);
	end component soc_video_system_video_decoder_0;

	component soc_video_system_video_dma_controller is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			stream_data          : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_startofpacket : in  std_logic                     := 'X';             -- startofpacket
			stream_endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			stream_valid         : in  std_logic                     := 'X';             -- valid
			stream_ready         : out std_logic;                                        -- ready
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_write         : out std_logic;                                        -- write
			master_writedata     : out std_logic_vector(7 downto 0)                      -- writedata
		);
	end component soc_video_system_video_dma_controller;

	component soc_video_system_video_dual_clock_buffer is
		port (
			clk_stream_in            : in  std_logic                     := 'X';             -- clk
			reset_stream_in          : in  std_logic                     := 'X';             -- reset
			clk_stream_out           : in  std_logic                     := 'X';             -- clk
			reset_stream_out         : in  std_logic                     := 'X';             -- reset
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_data           : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component soc_video_system_video_dual_clock_buffer;

	component soc_video_system_video_pixel_buffer_dma is
		port (
			clk                  : in  std_logic                     := 'X';             -- clk
			reset                : in  std_logic                     := 'X';             -- reset
			master_readdatavalid : in  std_logic                     := 'X';             -- readdatavalid
			master_waitrequest   : in  std_logic                     := 'X';             -- waitrequest
			master_address       : out std_logic_vector(31 downto 0);                    -- address
			master_arbiterlock   : out std_logic;                                        -- lock
			master_read          : out std_logic;                                        -- read
			master_readdata      : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			slave_address        : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			slave_byteenable     : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			slave_read           : in  std_logic                     := 'X';             -- read
			slave_write          : in  std_logic                     := 'X';             -- write
			slave_writedata      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			slave_readdata       : out std_logic_vector(31 downto 0);                    -- readdata
			stream_ready         : in  std_logic                     := 'X';             -- ready
			stream_startofpacket : out std_logic;                                        -- startofpacket
			stream_endofpacket   : out std_logic;                                        -- endofpacket
			stream_valid         : out std_logic;                                        -- valid
			stream_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component soc_video_system_video_pixel_buffer_dma;

	component soc_video_system_video_pixel_rgb_resampler_1 is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(29 downto 0)                     -- data
		);
	end component soc_video_system_video_pixel_rgb_resampler_1;

	component soc_video_system_video_pll is
		port (
			ref_clk_clk        : in  std_logic := 'X'; -- clk
			ref_reset_reset    : in  std_logic := 'X'; -- reset
			video_in_clk_clk   : out std_logic;        -- clk
			vga_clk_clk        : out std_logic;        -- clk
			reset_source_reset : out std_logic         -- reset
		);
	end component soc_video_system_video_pll;

	component soc_video_system_video_rgb_resampler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(7 downto 0)                      -- data
		);
	end component soc_video_system_video_rgb_resampler;

	component soc_video_system_video_scaler is
		port (
			clk                      : in  std_logic                     := 'X';             -- clk
			reset                    : in  std_logic                     := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                     := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                     := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                     := 'X';             -- valid
			stream_in_ready          : out std_logic;                                        -- ready
			stream_in_data           : in  std_logic_vector(23 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                     := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                        -- startofpacket
			stream_out_endofpacket   : out std_logic;                                        -- endofpacket
			stream_out_valid         : out std_logic;                                        -- valid
			stream_out_data          : out std_logic_vector(23 downto 0)                     -- data
		);
	end component soc_video_system_video_scaler;

	component soc_video_system_video_scaler_0 is
		port (
			clk                      : in  std_logic                    := 'X';             -- clk
			reset                    : in  std_logic                    := 'X';             -- reset
			stream_in_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid          : in  std_logic                    := 'X';             -- valid
			stream_in_ready          : out std_logic;                                       -- ready
			stream_in_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_out_ready         : in  std_logic                    := 'X';             -- ready
			stream_out_startofpacket : out std_logic;                                       -- startofpacket
			stream_out_endofpacket   : out std_logic;                                       -- endofpacket
			stream_out_valid         : out std_logic;                                       -- valid
			stream_out_data          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_channel       : out std_logic_vector(1 downto 0)                     -- channel
		);
	end component soc_video_system_video_scaler_0;

	component soc_video_system_video_stream_router_0 is
		port (
			clk                        : in  std_logic                    := 'X';             -- clk
			reset                      : in  std_logic                    := 'X';             -- reset
			stream_in_data             : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket    : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket      : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid            : in  std_logic                    := 'X';             -- valid
			stream_in_ready            : out std_logic;                                       -- ready
			stream_out_ready_0         : in  std_logic                    := 'X';             -- ready
			stream_out_data_0          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_startofpacket_0 : out std_logic;                                       -- startofpacket
			stream_out_endofpacket_0   : out std_logic;                                       -- endofpacket
			stream_out_valid_0         : out std_logic;                                       -- valid
			stream_out_ready_1         : in  std_logic                    := 'X';             -- ready
			stream_out_data_1          : out std_logic_vector(7 downto 0);                    -- data
			stream_out_startofpacket_1 : out std_logic;                                       -- startofpacket
			stream_out_endofpacket_1   : out std_logic;                                       -- endofpacket
			stream_out_valid_1         : out std_logic;                                       -- valid
			stream_select              : in  std_logic                    := 'X'              -- export
		);
	end component soc_video_system_video_stream_router_0;

	component soc_video_system_video_stream_router_1 is
		port (
			clk                       : in  std_logic                    := 'X';             -- clk
			reset                     : in  std_logic                    := 'X';             -- reset
			stream_in_data_0          : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket_0 : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket_0   : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid_0         : in  std_logic                    := 'X';             -- valid
			stream_in_ready_0         : out std_logic;                                       -- ready
			stream_in_data_1          : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			stream_in_startofpacket_1 : in  std_logic                    := 'X';             -- startofpacket
			stream_in_endofpacket_1   : in  std_logic                    := 'X';             -- endofpacket
			stream_in_valid_1         : in  std_logic                    := 'X';             -- valid
			stream_in_ready_1         : out std_logic;                                       -- ready
			stream_select             : in  std_logic                    := 'X';             -- export
			stream_out_ready          : in  std_logic                    := 'X';             -- ready
			stream_out_data           : out std_logic_vector(7 downto 0);                    -- data
			stream_out_startofpacket  : out std_logic;                                       -- startofpacket
			stream_out_endofpacket    : out std_logic;                                       -- endofpacket
			stream_out_valid          : out std_logic                                        -- valid
		);
	end component soc_video_system_video_stream_router_1;

	component soc_video_system_video_vga_controller is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset         : in  std_logic                     := 'X';             -- reset
			data          : in  std_logic_vector(29 downto 0) := (others => 'X'); -- data
			startofpacket : in  std_logic                     := 'X';             -- startofpacket
			endofpacket   : in  std_logic                     := 'X';             -- endofpacket
			valid         : in  std_logic                     := 'X';             -- valid
			ready         : out std_logic;                                        -- ready
			VGA_CLK       : out std_logic;                                        -- export
			VGA_HS        : out std_logic;                                        -- export
			VGA_VS        : out std_logic;                                        -- export
			VGA_BLANK     : out std_logic;                                        -- export
			VGA_SYNC      : out std_logic;                                        -- export
			VGA_R         : out std_logic_vector(7 downto 0);                     -- export
			VGA_G         : out std_logic_vector(7 downto 0);                     -- export
			VGA_B         : out std_logic_vector(7 downto 0)                      -- export
		);
	end component soc_video_system_video_vga_controller;

	component soc_video_system_mm_interconnect_0 is
		port (
			altpll_0_c0_clk                                              : in  std_logic                     := 'X';             -- clk
			clk_0_clk_clk                                                : in  std_logic                     := 'X';             -- clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset   : in  std_logic                     := 'X';             -- reset
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			video_dma_controller_reset_reset_bridge_in_reset_reset       : in  std_logic                     := 'X';             -- reset
			fpga_only_master_master_address                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			fpga_only_master_master_waitrequest                          : out std_logic;                                        -- waitrequest
			fpga_only_master_master_byteenable                           : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			fpga_only_master_master_read                                 : in  std_logic                     := 'X';             -- read
			fpga_only_master_master_readdata                             : out std_logic_vector(31 downto 0);                    -- readdata
			fpga_only_master_master_readdatavalid                        : out std_logic;                                        -- readdatavalid
			fpga_only_master_master_write                                : in  std_logic                     := 'X';             -- write
			fpga_only_master_master_writedata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			video_dma_controller_avalon_dma_master_address               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			video_dma_controller_avalon_dma_master_waitrequest           : out std_logic;                                        -- waitrequest
			video_dma_controller_avalon_dma_master_write                 : in  std_logic                     := 'X';             -- write
			video_dma_controller_avalon_dma_master_writedata             : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- writedata
			video_pixel_buffer_dma_avalon_pixel_dma_master_address       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- address
			video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest   : out std_logic;                                        -- waitrequest
			video_pixel_buffer_dma_avalon_pixel_dma_master_read          : in  std_logic                     := 'X';             -- read
			video_pixel_buffer_dma_avalon_pixel_dma_master_readdata      : out std_logic_vector(7 downto 0);                     -- readdata
			video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid : out std_logic;                                        -- readdatavalid
			video_pixel_buffer_dma_avalon_pixel_dma_master_lock          : in  std_logic                     := 'X';             -- lock
			altpll_0_pll_slave_address                                   : out std_logic_vector(1 downto 0);                     -- address
			altpll_0_pll_slave_write                                     : out std_logic;                                        -- write
			altpll_0_pll_slave_read                                      : out std_logic;                                        -- read
			altpll_0_pll_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			altpll_0_pll_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_address      : out std_logic_vector(1 downto 0);                     -- address
			audio_and_video_config_0_avalon_av_config_slave_write        : out std_logic;                                        -- write
			audio_and_video_config_0_avalon_av_config_slave_read         : out std_logic;                                        -- read
			audio_and_video_config_0_avalon_av_config_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata    : out std_logic_vector(31 downto 0);                    -- writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable   : out std_logic_vector(3 downto 0);                     -- byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest  : in  std_logic                     := 'X';             -- waitrequest
			pixel_buffer_s1_address                                      : out std_logic_vector(24 downto 0);                    -- address
			pixel_buffer_s1_write                                        : out std_logic;                                        -- write
			pixel_buffer_s1_read                                         : out std_logic;                                        -- read
			pixel_buffer_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			pixel_buffer_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			pixel_buffer_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			pixel_buffer_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			pixel_buffer_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			pixel_buffer_s1_chipselect                                   : out std_logic;                                        -- chipselect
			pixel_onchip_buffer_s1_address                               : out std_logic_vector(17 downto 0);                    -- address
			pixel_onchip_buffer_s1_write                                 : out std_logic;                                        -- write
			pixel_onchip_buffer_s1_readdata                              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			pixel_onchip_buffer_s1_writedata                             : out std_logic_vector(7 downto 0);                     -- writedata
			pixel_onchip_buffer_s1_chipselect                            : out std_logic;                                        -- chipselect
			pixel_onchip_buffer_s1_clken                                 : out std_logic;                                        -- clken
			video_dma_controller_avalon_dma_control_slave_address        : out std_logic_vector(1 downto 0);                     -- address
			video_dma_controller_avalon_dma_control_slave_write          : out std_logic;                                        -- write
			video_dma_controller_avalon_dma_control_slave_read           : out std_logic;                                        -- read
			video_dma_controller_avalon_dma_control_slave_readdata       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_dma_controller_avalon_dma_control_slave_writedata      : out std_logic_vector(31 downto 0);                    -- writedata
			video_dma_controller_avalon_dma_control_slave_byteenable     : out std_logic_vector(3 downto 0);                     -- byteenable
			video_pixel_buffer_dma_avalon_control_slave_address          : out std_logic_vector(1 downto 0);                     -- address
			video_pixel_buffer_dma_avalon_control_slave_write            : out std_logic;                                        -- write
			video_pixel_buffer_dma_avalon_control_slave_read             : out std_logic;                                        -- read
			video_pixel_buffer_dma_avalon_control_slave_readdata         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			video_pixel_buffer_dma_avalon_control_slave_writedata        : out std_logic_vector(31 downto 0);                    -- writedata
			video_pixel_buffer_dma_avalon_control_slave_byteenable       : out std_logic_vector(3 downto 0)                      -- byteenable
		);
	end component soc_video_system_mm_interconnect_0;

	component soc_video_system_avalon_st_adapter is
		generic (
			inBitsPerSymbol : integer := 8;
			inUsePackets    : integer := 0;
			inDataWidth     : integer := 8;
			inChannelWidth  : integer := 3;
			inErrorWidth    : integer := 2;
			inUseEmptyPort  : integer := 0;
			inUseValid      : integer := 1;
			inUseReady      : integer := 1;
			inReadyLatency  : integer := 0;
			outDataWidth    : integer := 32;
			outChannelWidth : integer := 3;
			outErrorWidth   : integer := 2;
			outUseEmptyPort : integer := 0;
			outUseValid     : integer := 1;
			outUseReady     : integer := 1;
			outReadyLatency : integer := 0
		);
		port (
			in_clk_0_clk        : in  std_logic                    := 'X';             -- clk
			in_rst_0_reset      : in  std_logic                    := 'X';             -- reset
			in_0_data           : in  std_logic_vector(7 downto 0) := (others => 'X'); -- data
			in_0_valid          : in  std_logic                    := 'X';             -- valid
			in_0_ready          : out std_logic;                                       -- ready
			in_0_startofpacket  : in  std_logic                    := 'X';             -- startofpacket
			in_0_endofpacket    : in  std_logic                    := 'X';             -- endofpacket
			in_0_channel        : in  std_logic_vector(1 downto 0) := (others => 'X'); -- channel
			out_0_data          : out std_logic_vector(7 downto 0);                    -- data
			out_0_valid         : out std_logic;                                       -- valid
			out_0_ready         : in  std_logic                    := 'X';             -- ready
			out_0_startofpacket : out std_logic;                                       -- startofpacket
			out_0_endofpacket   : out std_logic                                        -- endofpacket
		);
	end component soc_video_system_avalon_st_adapter;

	component altera_reset_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_in2      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component altera_reset_controller;

	signal video_bayer_resampler_avalon_bayer_source_valid                               : std_logic;                     -- video_bayer_resampler:stream_out_valid -> video_clipper:stream_in_valid
	signal video_bayer_resampler_avalon_bayer_source_data                                : std_logic_vector(23 downto 0); -- video_bayer_resampler:stream_out_data -> video_clipper:stream_in_data
	signal video_bayer_resampler_avalon_bayer_source_ready                               : std_logic;                     -- video_clipper:stream_in_ready -> video_bayer_resampler:stream_out_ready
	signal video_bayer_resampler_avalon_bayer_source_startofpacket                       : std_logic;                     -- video_bayer_resampler:stream_out_startofpacket -> video_clipper:stream_in_startofpacket
	signal video_bayer_resampler_avalon_bayer_source_endofpacket                         : std_logic;                     -- video_bayer_resampler:stream_out_endofpacket -> video_clipper:stream_in_endofpacket
	signal video_clipper_avalon_clipper_source_valid                                     : std_logic;                     -- video_clipper:stream_out_valid -> video_scaler:stream_in_valid
	signal video_clipper_avalon_clipper_source_data                                      : std_logic_vector(23 downto 0); -- video_clipper:stream_out_data -> video_scaler:stream_in_data
	signal video_clipper_avalon_clipper_source_ready                                     : std_logic;                     -- video_scaler:stream_in_ready -> video_clipper:stream_out_ready
	signal video_clipper_avalon_clipper_source_startofpacket                             : std_logic;                     -- video_clipper:stream_out_startofpacket -> video_scaler:stream_in_startofpacket
	signal video_clipper_avalon_clipper_source_endofpacket                               : std_logic;                     -- video_clipper:stream_out_endofpacket -> video_scaler:stream_in_endofpacket
	signal video_dual_clock_buffer_avalon_dc_buffer_source_valid                         : std_logic;                     -- video_dual_clock_buffer:stream_out_valid -> video_vga_controller:valid
	signal video_dual_clock_buffer_avalon_dc_buffer_source_data                          : std_logic_vector(29 downto 0); -- video_dual_clock_buffer:stream_out_data -> video_vga_controller:data
	signal video_dual_clock_buffer_avalon_dc_buffer_source_ready                         : std_logic;                     -- video_vga_controller:ready -> video_dual_clock_buffer:stream_out_ready
	signal video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket                 : std_logic;                     -- video_dual_clock_buffer:stream_out_startofpacket -> video_vga_controller:startofpacket
	signal video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket                   : std_logic;                     -- video_dual_clock_buffer:stream_out_endofpacket -> video_vga_controller:endofpacket
	signal video_decoder_0_avalon_decoder_source_valid                                   : std_logic;                     -- video_decoder_0:stream_out_valid -> video_bayer_resampler:stream_in_valid
	signal video_decoder_0_avalon_decoder_source_data                                    : std_logic_vector(7 downto 0);  -- video_decoder_0:stream_out_data -> video_bayer_resampler:stream_in_data
	signal video_decoder_0_avalon_decoder_source_ready                                   : std_logic;                     -- video_bayer_resampler:stream_in_ready -> video_decoder_0:stream_out_ready
	signal video_decoder_0_avalon_decoder_source_startofpacket                           : std_logic;                     -- video_decoder_0:stream_out_startofpacket -> video_bayer_resampler:stream_in_startofpacket
	signal video_decoder_0_avalon_decoder_source_endofpacket                             : std_logic;                     -- video_decoder_0:stream_out_endofpacket -> video_bayer_resampler:stream_in_endofpacket
	signal video_pixel_buffer_dma_avalon_pixel_source_valid                              : std_logic;                     -- video_pixel_buffer_dma:stream_valid -> video_scaler_0:stream_in_valid
	signal video_pixel_buffer_dma_avalon_pixel_source_data                               : std_logic_vector(7 downto 0);  -- video_pixel_buffer_dma:stream_data -> video_scaler_0:stream_in_data
	signal video_pixel_buffer_dma_avalon_pixel_source_ready                              : std_logic;                     -- video_scaler_0:stream_in_ready -> video_pixel_buffer_dma:stream_ready
	signal video_pixel_buffer_dma_avalon_pixel_source_startofpacket                      : std_logic;                     -- video_pixel_buffer_dma:stream_startofpacket -> video_scaler_0:stream_in_startofpacket
	signal video_pixel_buffer_dma_avalon_pixel_source_endofpacket                        : std_logic;                     -- video_pixel_buffer_dma:stream_endofpacket -> video_scaler_0:stream_in_endofpacket
	signal video_pixel_rgb_resampler_1_avalon_rgb_source_valid                           : std_logic;                     -- video_pixel_rgb_resampler_1:stream_out_valid -> video_dual_clock_buffer:stream_in_valid
	signal video_pixel_rgb_resampler_1_avalon_rgb_source_data                            : std_logic_vector(29 downto 0); -- video_pixel_rgb_resampler_1:stream_out_data -> video_dual_clock_buffer:stream_in_data
	signal video_pixel_rgb_resampler_1_avalon_rgb_source_ready                           : std_logic;                     -- video_dual_clock_buffer:stream_in_ready -> video_pixel_rgb_resampler_1:stream_out_ready
	signal video_pixel_rgb_resampler_1_avalon_rgb_source_startofpacket                   : std_logic;                     -- video_pixel_rgb_resampler_1:stream_out_startofpacket -> video_dual_clock_buffer:stream_in_startofpacket
	signal video_pixel_rgb_resampler_1_avalon_rgb_source_endofpacket                     : std_logic;                     -- video_pixel_rgb_resampler_1:stream_out_endofpacket -> video_dual_clock_buffer:stream_in_endofpacket
	signal video_rgb_resampler_avalon_rgb_source_valid                                   : std_logic;                     -- video_rgb_resampler:stream_out_valid -> video_stream_router_0:stream_in_valid
	signal video_rgb_resampler_avalon_rgb_source_data                                    : std_logic_vector(7 downto 0);  -- video_rgb_resampler:stream_out_data -> video_stream_router_0:stream_in_data
	signal video_rgb_resampler_avalon_rgb_source_ready                                   : std_logic;                     -- video_stream_router_0:stream_in_ready -> video_rgb_resampler:stream_out_ready
	signal video_rgb_resampler_avalon_rgb_source_startofpacket                           : std_logic;                     -- video_rgb_resampler:stream_out_startofpacket -> video_stream_router_0:stream_in_startofpacket
	signal video_rgb_resampler_avalon_rgb_source_endofpacket                             : std_logic;                     -- video_rgb_resampler:stream_out_endofpacket -> video_stream_router_0:stream_in_endofpacket
	signal video_scaler_avalon_scaler_source_valid                                       : std_logic;                     -- video_scaler:stream_out_valid -> video_rgb_resampler:stream_in_valid
	signal video_scaler_avalon_scaler_source_data                                        : std_logic_vector(23 downto 0); -- video_scaler:stream_out_data -> video_rgb_resampler:stream_in_data
	signal video_scaler_avalon_scaler_source_ready                                       : std_logic;                     -- video_rgb_resampler:stream_in_ready -> video_scaler:stream_out_ready
	signal video_scaler_avalon_scaler_source_startofpacket                               : std_logic;                     -- video_scaler:stream_out_startofpacket -> video_rgb_resampler:stream_in_startofpacket
	signal video_scaler_avalon_scaler_source_endofpacket                                 : std_logic;                     -- video_scaler:stream_out_endofpacket -> video_rgb_resampler:stream_in_endofpacket
	signal video_stream_router_1_avalon_stream_router_source_valid                       : std_logic;                     -- video_stream_router_1:stream_out_valid -> video_dma_controller:stream_valid
	signal video_stream_router_1_avalon_stream_router_source_data                        : std_logic_vector(7 downto 0);  -- video_stream_router_1:stream_out_data -> video_dma_controller:stream_data
	signal video_stream_router_1_avalon_stream_router_source_ready                       : std_logic;                     -- video_dma_controller:stream_ready -> video_stream_router_1:stream_out_ready
	signal video_stream_router_1_avalon_stream_router_source_startofpacket               : std_logic;                     -- video_stream_router_1:stream_out_startofpacket -> video_dma_controller:stream_startofpacket
	signal video_stream_router_1_avalon_stream_router_source_endofpacket                 : std_logic;                     -- video_stream_router_1:stream_out_endofpacket -> video_dma_controller:stream_endofpacket
	signal video_stream_router_0_avalon_stream_router_source_0_valid                     : std_logic;                     -- video_stream_router_0:stream_out_valid_0 -> video_stream_router_1:stream_in_valid_0
	signal video_stream_router_0_avalon_stream_router_source_0_data                      : std_logic_vector(7 downto 0);  -- video_stream_router_0:stream_out_data_0 -> video_stream_router_1:stream_in_data_0
	signal video_stream_router_0_avalon_stream_router_source_0_ready                     : std_logic;                     -- video_stream_router_1:stream_in_ready_0 -> video_stream_router_0:stream_out_ready_0
	signal video_stream_router_0_avalon_stream_router_source_0_startofpacket             : std_logic;                     -- video_stream_router_0:stream_out_startofpacket_0 -> video_stream_router_1:stream_in_startofpacket_0
	signal video_stream_router_0_avalon_stream_router_source_0_endofpacket               : std_logic;                     -- video_stream_router_0:stream_out_endofpacket_0 -> video_stream_router_1:stream_in_endofpacket_0
	signal video_stream_router_0_avalon_stream_router_source_1_valid                     : std_logic;                     -- video_stream_router_0:stream_out_valid_1 -> sobel_edge_detector_0:in_valid
	signal video_stream_router_0_avalon_stream_router_source_1_data                      : std_logic_vector(7 downto 0);  -- video_stream_router_0:stream_out_data_1 -> sobel_edge_detector_0:in_data
	signal video_stream_router_0_avalon_stream_router_source_1_ready                     : std_logic;                     -- sobel_edge_detector_0:in_ready -> video_stream_router_0:stream_out_ready_1
	signal video_stream_router_0_avalon_stream_router_source_1_startofpacket             : std_logic;                     -- video_stream_router_0:stream_out_startofpacket_1 -> sobel_edge_detector_0:in_startofpacket
	signal video_stream_router_0_avalon_stream_router_source_1_endofpacket               : std_logic;                     -- video_stream_router_0:stream_out_endofpacket_1 -> sobel_edge_detector_0:in_endofpacket
	signal sobel_edge_detector_0_avalon_streaming_source_valid                           : std_logic;                     -- sobel_edge_detector_0:out_valid -> video_stream_router_1:stream_in_valid_1
	signal sobel_edge_detector_0_avalon_streaming_source_data                            : std_logic_vector(7 downto 0);  -- sobel_edge_detector_0:out_data -> video_stream_router_1:stream_in_data_1
	signal sobel_edge_detector_0_avalon_streaming_source_ready                           : std_logic;                     -- video_stream_router_1:stream_in_ready_1 -> sobel_edge_detector_0:out_ready
	signal sobel_edge_detector_0_avalon_streaming_source_startofpacket                   : std_logic;                     -- sobel_edge_detector_0:out_startofpacket -> video_stream_router_1:stream_in_startofpacket_1
	signal sobel_edge_detector_0_avalon_streaming_source_endofpacket                     : std_logic;                     -- sobel_edge_detector_0:out_endofpacket -> video_stream_router_1:stream_in_endofpacket_1
	signal altpll_0_c0_clk                                                               : std_logic;                     -- altpll_0:c0 -> [audio_and_video_config_0:clk, avalon_st_adapter:in_clk_0_clk, fpga_only_master:clk_clk, mm_interconnect_0:altpll_0_c0_clk, pixel_buffer:clk, pixel_onchip_buffer:clk, rst_controller_001:clk, sobel_edge_detector_0:clk, video_bayer_resampler:clk, video_clipper:clk, video_decoder_0:clk, video_dma_controller:clk, video_dual_clock_buffer:clk_stream_in, video_pixel_buffer_dma:clk, video_pixel_rgb_resampler_1:clk, video_rgb_resampler:clk, video_scaler:clk, video_scaler_0:clk, video_stream_router_0:clk, video_stream_router_1:clk]
	signal video_pll_vga_clk_clk                                                         : std_logic;                     -- video_pll:vga_clk_clk -> [rst_controller_003:clk, video_dual_clock_buffer:clk_stream_out, video_vga_controller:clk]
	signal video_dma_controller_avalon_dma_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:video_dma_controller_avalon_dma_master_waitrequest -> video_dma_controller:master_waitrequest
	signal video_dma_controller_avalon_dma_master_address                                : std_logic_vector(31 downto 0); -- video_dma_controller:master_address -> mm_interconnect_0:video_dma_controller_avalon_dma_master_address
	signal video_dma_controller_avalon_dma_master_write                                  : std_logic;                     -- video_dma_controller:master_write -> mm_interconnect_0:video_dma_controller_avalon_dma_master_write
	signal video_dma_controller_avalon_dma_master_writedata                              : std_logic_vector(7 downto 0);  -- video_dma_controller:master_writedata -> mm_interconnect_0:video_dma_controller_avalon_dma_master_writedata
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest                    : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest -> video_pixel_buffer_dma:master_waitrequest
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_readdata                       : std_logic_vector(7 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_readdata -> video_pixel_buffer_dma:master_readdata
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_address                        : std_logic_vector(31 downto 0); -- video_pixel_buffer_dma:master_address -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_address
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_read                           : std_logic;                     -- video_pixel_buffer_dma:master_read -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_read
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid                  : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid -> video_pixel_buffer_dma:master_readdatavalid
	signal video_pixel_buffer_dma_avalon_pixel_dma_master_lock                           : std_logic;                     -- video_pixel_buffer_dma:master_arbiterlock -> mm_interconnect_0:video_pixel_buffer_dma_avalon_pixel_dma_master_lock
	signal fpga_only_master_master_readdata                                              : std_logic_vector(31 downto 0); -- mm_interconnect_0:fpga_only_master_master_readdata -> fpga_only_master:master_readdata
	signal fpga_only_master_master_waitrequest                                           : std_logic;                     -- mm_interconnect_0:fpga_only_master_master_waitrequest -> fpga_only_master:master_waitrequest
	signal fpga_only_master_master_address                                               : std_logic_vector(31 downto 0); -- fpga_only_master:master_address -> mm_interconnect_0:fpga_only_master_master_address
	signal fpga_only_master_master_read                                                  : std_logic;                     -- fpga_only_master:master_read -> mm_interconnect_0:fpga_only_master_master_read
	signal fpga_only_master_master_byteenable                                            : std_logic_vector(3 downto 0);  -- fpga_only_master:master_byteenable -> mm_interconnect_0:fpga_only_master_master_byteenable
	signal fpga_only_master_master_readdatavalid                                         : std_logic;                     -- mm_interconnect_0:fpga_only_master_master_readdatavalid -> fpga_only_master:master_readdatavalid
	signal fpga_only_master_master_write                                                 : std_logic;                     -- fpga_only_master:master_write -> mm_interconnect_0:fpga_only_master_master_write
	signal fpga_only_master_master_writedata                                             : std_logic_vector(31 downto 0); -- fpga_only_master:master_writedata -> mm_interconnect_0:fpga_only_master_master_writedata
	signal mm_interconnect_0_pixel_onchip_buffer_s1_chipselect                           : std_logic;                     -- mm_interconnect_0:pixel_onchip_buffer_s1_chipselect -> pixel_onchip_buffer:chipselect
	signal mm_interconnect_0_pixel_onchip_buffer_s1_readdata                             : std_logic_vector(7 downto 0);  -- pixel_onchip_buffer:readdata -> mm_interconnect_0:pixel_onchip_buffer_s1_readdata
	signal mm_interconnect_0_pixel_onchip_buffer_s1_address                              : std_logic_vector(17 downto 0); -- mm_interconnect_0:pixel_onchip_buffer_s1_address -> pixel_onchip_buffer:address
	signal mm_interconnect_0_pixel_onchip_buffer_s1_write                                : std_logic;                     -- mm_interconnect_0:pixel_onchip_buffer_s1_write -> pixel_onchip_buffer:write
	signal mm_interconnect_0_pixel_onchip_buffer_s1_writedata                            : std_logic_vector(7 downto 0);  -- mm_interconnect_0:pixel_onchip_buffer_s1_writedata -> pixel_onchip_buffer:writedata
	signal mm_interconnect_0_pixel_onchip_buffer_s1_clken                                : std_logic;                     -- mm_interconnect_0:pixel_onchip_buffer_s1_clken -> pixel_onchip_buffer:clken
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata    : std_logic_vector(31 downto 0); -- audio_and_video_config_0:readdata -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_readdata
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest : std_logic;                     -- audio_and_video_config_0:waitrequest -> mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_waitrequest
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address     : std_logic_vector(1 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_address -> audio_and_video_config_0:address
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read        : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_read -> audio_and_video_config_0:read
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable  : std_logic_vector(3 downto 0);  -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_byteenable -> audio_and_video_config_0:byteenable
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write       : std_logic;                     -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_write -> audio_and_video_config_0:write
	signal mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata   : std_logic_vector(31 downto 0); -- mm_interconnect_0:audio_and_video_config_0_avalon_av_config_slave_writedata -> audio_and_video_config_0:writedata
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata        : std_logic_vector(31 downto 0); -- video_pixel_buffer_dma:slave_readdata -> mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_readdata
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_address -> video_pixel_buffer_dma:slave_address
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read            : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_read -> video_pixel_buffer_dma:slave_read
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable      : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_byteenable -> video_pixel_buffer_dma:slave_byteenable
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write           : std_logic;                     -- mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_write -> video_pixel_buffer_dma:slave_write
	signal mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_pixel_buffer_dma_avalon_control_slave_writedata -> video_pixel_buffer_dma:slave_writedata
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_readdata      : std_logic_vector(31 downto 0); -- video_dma_controller:slave_readdata -> mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_readdata
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_address       : std_logic_vector(1 downto 0);  -- mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_address -> video_dma_controller:slave_address
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_read          : std_logic;                     -- mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_read -> video_dma_controller:slave_read
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_byteenable    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_byteenable -> video_dma_controller:slave_byteenable
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_write         : std_logic;                     -- mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_write -> video_dma_controller:slave_write
	signal mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_writedata     : std_logic_vector(31 downto 0); -- mm_interconnect_0:video_dma_controller_avalon_dma_control_slave_writedata -> video_dma_controller:slave_writedata
	signal mm_interconnect_0_altpll_0_pll_slave_readdata                                 : std_logic_vector(31 downto 0); -- altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	signal mm_interconnect_0_altpll_0_pll_slave_address                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	signal mm_interconnect_0_altpll_0_pll_slave_read                                     : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	signal mm_interconnect_0_altpll_0_pll_slave_write                                    : std_logic;                     -- mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	signal mm_interconnect_0_altpll_0_pll_slave_writedata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	signal mm_interconnect_0_pixel_buffer_s1_chipselect                                  : std_logic;                     -- mm_interconnect_0:pixel_buffer_s1_chipselect -> pixel_buffer:az_cs
	signal mm_interconnect_0_pixel_buffer_s1_readdata                                    : std_logic_vector(15 downto 0); -- pixel_buffer:za_data -> mm_interconnect_0:pixel_buffer_s1_readdata
	signal mm_interconnect_0_pixel_buffer_s1_waitrequest                                 : std_logic;                     -- pixel_buffer:za_waitrequest -> mm_interconnect_0:pixel_buffer_s1_waitrequest
	signal mm_interconnect_0_pixel_buffer_s1_address                                     : std_logic_vector(24 downto 0); -- mm_interconnect_0:pixel_buffer_s1_address -> pixel_buffer:az_addr
	signal mm_interconnect_0_pixel_buffer_s1_read                                        : std_logic;                     -- mm_interconnect_0:pixel_buffer_s1_read -> mm_interconnect_0_pixel_buffer_s1_read:in
	signal mm_interconnect_0_pixel_buffer_s1_byteenable                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pixel_buffer_s1_byteenable -> mm_interconnect_0_pixel_buffer_s1_byteenable:in
	signal mm_interconnect_0_pixel_buffer_s1_readdatavalid                               : std_logic;                     -- pixel_buffer:za_valid -> mm_interconnect_0:pixel_buffer_s1_readdatavalid
	signal mm_interconnect_0_pixel_buffer_s1_write                                       : std_logic;                     -- mm_interconnect_0:pixel_buffer_s1_write -> mm_interconnect_0_pixel_buffer_s1_write:in
	signal mm_interconnect_0_pixel_buffer_s1_writedata                                   : std_logic_vector(15 downto 0); -- mm_interconnect_0:pixel_buffer_s1_writedata -> pixel_buffer:az_data
	signal video_scaler_0_avalon_scaler_source_valid                                     : std_logic;                     -- video_scaler_0:stream_out_valid -> avalon_st_adapter:in_0_valid
	signal video_scaler_0_avalon_scaler_source_data                                      : std_logic_vector(7 downto 0);  -- video_scaler_0:stream_out_data -> avalon_st_adapter:in_0_data
	signal video_scaler_0_avalon_scaler_source_ready                                     : std_logic;                     -- avalon_st_adapter:in_0_ready -> video_scaler_0:stream_out_ready
	signal video_scaler_0_avalon_scaler_source_channel                                   : std_logic_vector(1 downto 0);  -- video_scaler_0:stream_out_channel -> avalon_st_adapter:in_0_channel
	signal video_scaler_0_avalon_scaler_source_startofpacket                             : std_logic;                     -- video_scaler_0:stream_out_startofpacket -> avalon_st_adapter:in_0_startofpacket
	signal video_scaler_0_avalon_scaler_source_endofpacket                               : std_logic;                     -- video_scaler_0:stream_out_endofpacket -> avalon_st_adapter:in_0_endofpacket
	signal avalon_st_adapter_out_0_valid                                                 : std_logic;                     -- avalon_st_adapter:out_0_valid -> video_pixel_rgb_resampler_1:stream_in_valid
	signal avalon_st_adapter_out_0_data                                                  : std_logic_vector(7 downto 0);  -- avalon_st_adapter:out_0_data -> video_pixel_rgb_resampler_1:stream_in_data
	signal avalon_st_adapter_out_0_ready                                                 : std_logic;                     -- video_pixel_rgb_resampler_1:stream_in_ready -> avalon_st_adapter:out_0_ready
	signal avalon_st_adapter_out_0_startofpacket                                         : std_logic;                     -- avalon_st_adapter:out_0_startofpacket -> video_pixel_rgb_resampler_1:stream_in_startofpacket
	signal avalon_st_adapter_out_0_endofpacket                                           : std_logic;                     -- avalon_st_adapter:out_0_endofpacket -> video_pixel_rgb_resampler_1:stream_in_endofpacket
	signal rst_controller_reset_out_reset                                                : std_logic;                     -- rst_controller:reset_out -> [altpll_0:reset, mm_interconnect_0:altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset, video_pll:ref_reset_reset]
	signal fpga_only_master_master_reset_reset                                           : std_logic;                     -- fpga_only_master:master_reset_reset -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	signal video_pll_reset_source_reset                                                  : std_logic;                     -- video_pll:reset_source_reset -> [rst_controller:reset_in2, rst_controller_001:reset_in2, rst_controller_002:reset_in2, rst_controller_003:reset_in2]
	signal rst_controller_001_reset_out_reset                                            : std_logic;                     -- rst_controller_001:reset_out -> [audio_and_video_config_0:reset, avalon_st_adapter:in_rst_0_reset, mm_interconnect_0:fpga_only_master_clk_reset_reset_bridge_in_reset_reset, mm_interconnect_0:video_dma_controller_reset_reset_bridge_in_reset_reset, pixel_onchip_buffer:reset, rst_controller_001_reset_out_reset:in, sobel_edge_detector_0:reset, video_bayer_resampler:reset, video_clipper:reset, video_decoder_0:reset, video_dma_controller:reset, video_dual_clock_buffer:reset_stream_in, video_pixel_buffer_dma:reset, video_pixel_rgb_resampler_1:reset, video_rgb_resampler:reset, video_scaler:reset, video_scaler_0:reset, video_stream_router_0:reset, video_stream_router_1:reset]
	signal rst_controller_002_reset_out_reset                                            : std_logic;                     -- rst_controller_002:reset_out -> fpga_only_master:clk_reset_reset
	signal rst_controller_003_reset_out_reset                                            : std_logic;                     -- rst_controller_003:reset_out -> [video_dual_clock_buffer:reset_stream_out, video_vga_controller:reset]
	signal reset_reset_n_ports_inv                                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_pixel_buffer_s1_read_ports_inv                              : std_logic;                     -- mm_interconnect_0_pixel_buffer_s1_read:inv -> pixel_buffer:az_rd_n
	signal mm_interconnect_0_pixel_buffer_s1_byteenable_ports_inv                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0_pixel_buffer_s1_byteenable:inv -> pixel_buffer:az_be_n
	signal mm_interconnect_0_pixel_buffer_s1_write_ports_inv                             : std_logic;                     -- mm_interconnect_0_pixel_buffer_s1_write:inv -> pixel_buffer:az_wr_n
	signal rst_controller_001_reset_out_reset_ports_inv                                  : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> pixel_buffer:reset_n

begin

	altpll_0 : component soc_video_system_altpll_0
		port map (
			clk                => clk_clk,                                        --       inclk_interface.clk
			reset              => rst_controller_reset_out_reset,                 -- inclk_interface_reset.reset
			read               => mm_interconnect_0_altpll_0_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_altpll_0_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_altpll_0_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_altpll_0_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_altpll_0_pll_slave_writedata, --                      .writedata
			c0                 => altpll_0_c0_clk,                                --                    c0.clk
			c1                 => clk_sdram_clk,                                  --                    c1.clk
			scandone           => open,                                           --           (terminated)
			scandataout        => open,                                           --           (terminated)
			c2                 => open,                                           --           (terminated)
			c3                 => open,                                           --           (terminated)
			c4                 => open,                                           --           (terminated)
			areset             => '0',                                            --           (terminated)
			locked             => open,                                           --           (terminated)
			phasedone          => open,                                           --           (terminated)
			phasecounterselect => "000",                                          --           (terminated)
			phaseupdown        => '0',                                            --           (terminated)
			phasestep          => '0',                                            --           (terminated)
			scanclk            => '0',                                            --           (terminated)
			scanclkena         => '0',                                            --           (terminated)
			scandata           => '0',                                            --           (terminated)
			configupdate       => '0'                                             --           (terminated)
		);

	audio_and_video_config_0 : component soc_video_system_audio_and_video_config_0
		port map (
			clk         => altpll_0_c0_clk,                                                               --                    clk.clk
			reset       => rst_controller_001_reset_out_reset,                                            --                  reset.reset
			address     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     -- avalon_av_config_slave.address
			byteenable  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                       .byteenable
			read        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                       .read
			write       => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                       .write
			writedata   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                       .writedata
			readdata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                       .readdata
			waitrequest => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                       .waitrequest
			I2C_SDAT    => video_config_SDAT,                                                             --     external_interface.export
			I2C_SCLK    => video_config_SCLK                                                              --                       .export
		);

	fpga_only_master : component soc_video_system_fpga_only_master
		generic map (
			USE_PLI     => 0,
			PLI_PORT    => 50000,
			FIFO_DEPTHS => 2
		)
		port map (
			clk_clk              => altpll_0_c0_clk,                       --          clk.clk
			clk_reset_reset      => rst_controller_002_reset_out_reset,    --    clk_reset.reset
			master_address       => fpga_only_master_master_address,       --       master.address
			master_readdata      => fpga_only_master_master_readdata,      --             .readdata
			master_read          => fpga_only_master_master_read,          --             .read
			master_write         => fpga_only_master_master_write,         --             .write
			master_writedata     => fpga_only_master_master_writedata,     --             .writedata
			master_waitrequest   => fpga_only_master_master_waitrequest,   --             .waitrequest
			master_readdatavalid => fpga_only_master_master_readdatavalid, --             .readdatavalid
			master_byteenable    => fpga_only_master_master_byteenable,    --             .byteenable
			master_reset_reset   => fpga_only_master_master_reset_reset    -- master_reset.reset
		);

	pixel_buffer : component soc_video_system_pixel_buffer
		port map (
			clk            => altpll_0_c0_clk,                                        --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,           -- reset.reset_n
			az_addr        => mm_interconnect_0_pixel_buffer_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_pixel_buffer_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_pixel_buffer_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_pixel_buffer_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_pixel_buffer_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_pixel_buffer_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_pixel_buffer_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_pixel_buffer_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_pixel_buffer_s1_waitrequest,          --      .waitrequest
			zs_addr        => video_sdram_addr,                                       --  wire.export
			zs_ba          => video_sdram_ba,                                         --      .export
			zs_cas_n       => video_sdram_cas_n,                                      --      .export
			zs_cke         => video_sdram_cke,                                        --      .export
			zs_cs_n        => video_sdram_cs_n,                                       --      .export
			zs_dq          => video_sdram_dq,                                         --      .export
			zs_dqm         => video_sdram_dqm,                                        --      .export
			zs_ras_n       => video_sdram_ras_n,                                      --      .export
			zs_we_n        => video_sdram_we_n                                        --      .export
		);

	pixel_onchip_buffer : component soc_video_system_pixel_onchip_buffer
		port map (
			clk        => altpll_0_c0_clk,                                     --   clk1.clk
			address    => mm_interconnect_0_pixel_onchip_buffer_s1_address,    --     s1.address
			clken      => mm_interconnect_0_pixel_onchip_buffer_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_pixel_onchip_buffer_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_pixel_onchip_buffer_s1_write,      --       .write
			readdata   => mm_interconnect_0_pixel_onchip_buffer_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_pixel_onchip_buffer_s1_writedata,  --       .writedata
			reset      => rst_controller_001_reset_out_reset,                  -- reset1.reset
			reset_req  => '0',                                                 -- (terminated)
			freeze     => '0'                                                  -- (terminated)
		);

	sobel_edge_detector_0 : component altera_up_avalon_video_edge_detection
		generic map (
			WIDTH => 320
		)
		port map (
			clk               => altpll_0_c0_clk,                                                   --                   clock.clk
			reset             => rst_controller_001_reset_out_reset,                                --                   reset.reset
			bypass            => edge_detect_bypass,                                                --             conduit_end.bypass
			in_data           => video_stream_router_0_avalon_stream_router_source_1_data,          --   avalon_streaming_sink.data
			in_startofpacket  => video_stream_router_0_avalon_stream_router_source_1_startofpacket, --                        .startofpacket
			in_endofpacket    => video_stream_router_0_avalon_stream_router_source_1_endofpacket,   --                        .endofpacket
			in_valid          => video_stream_router_0_avalon_stream_router_source_1_valid,         --                        .valid
			in_ready          => video_stream_router_0_avalon_stream_router_source_1_ready,         --                        .ready
			out_data          => sobel_edge_detector_0_avalon_streaming_source_data,                -- avalon_streaming_source.data
			out_startofpacket => sobel_edge_detector_0_avalon_streaming_source_startofpacket,       --                        .startofpacket
			out_endofpacket   => sobel_edge_detector_0_avalon_streaming_source_endofpacket,         --                        .endofpacket
			out_valid         => sobel_edge_detector_0_avalon_streaming_source_valid,               --                        .valid
			out_ready         => sobel_edge_detector_0_avalon_streaming_source_ready                --                        .ready
		);

	video_bayer_resampler : component soc_video_system_video_bayer_resampler
		port map (
			clk                      => altpll_0_c0_clk,                                         --                 clk.clk
			reset                    => rst_controller_001_reset_out_reset,                      --               reset.reset
			stream_in_data           => video_decoder_0_avalon_decoder_source_data,              --   avalon_bayer_sink.data
			stream_in_startofpacket  => video_decoder_0_avalon_decoder_source_startofpacket,     --                    .startofpacket
			stream_in_endofpacket    => video_decoder_0_avalon_decoder_source_endofpacket,       --                    .endofpacket
			stream_in_valid          => video_decoder_0_avalon_decoder_source_valid,             --                    .valid
			stream_in_ready          => video_decoder_0_avalon_decoder_source_ready,             --                    .ready
			stream_out_ready         => video_bayer_resampler_avalon_bayer_source_ready,         -- avalon_bayer_source.ready
			stream_out_data          => video_bayer_resampler_avalon_bayer_source_data,          --                    .data
			stream_out_startofpacket => video_bayer_resampler_avalon_bayer_source_startofpacket, --                    .startofpacket
			stream_out_endofpacket   => video_bayer_resampler_avalon_bayer_source_endofpacket,   --                    .endofpacket
			stream_out_valid         => video_bayer_resampler_avalon_bayer_source_valid          --                    .valid
		);

	video_clipper : component soc_video_system_video_clipper
		port map (
			clk                      => altpll_0_c0_clk,                                         --                   clk.clk
			reset                    => rst_controller_001_reset_out_reset,                      --                 reset.reset
			stream_in_data           => video_bayer_resampler_avalon_bayer_source_data,          --   avalon_clipper_sink.data
			stream_in_startofpacket  => video_bayer_resampler_avalon_bayer_source_startofpacket, --                      .startofpacket
			stream_in_endofpacket    => video_bayer_resampler_avalon_bayer_source_endofpacket,   --                      .endofpacket
			stream_in_valid          => video_bayer_resampler_avalon_bayer_source_valid,         --                      .valid
			stream_in_ready          => video_bayer_resampler_avalon_bayer_source_ready,         --                      .ready
			stream_out_ready         => video_clipper_avalon_clipper_source_ready,               -- avalon_clipper_source.ready
			stream_out_data          => video_clipper_avalon_clipper_source_data,                --                      .data
			stream_out_startofpacket => video_clipper_avalon_clipper_source_startofpacket,       --                      .startofpacket
			stream_out_endofpacket   => video_clipper_avalon_clipper_source_endofpacket,         --                      .endofpacket
			stream_out_valid         => video_clipper_avalon_clipper_source_valid                --                      .valid
		);

	video_decoder_0 : component soc_video_system_video_decoder_0
		port map (
			clk                      => altpll_0_c0_clk,                                     --                   clk.clk
			reset                    => rst_controller_001_reset_out_reset,                  --                 reset.reset
			stream_out_ready         => video_decoder_0_avalon_decoder_source_ready,         -- avalon_decoder_source.ready
			stream_out_startofpacket => video_decoder_0_avalon_decoder_source_startofpacket, --                      .startofpacket
			stream_out_endofpacket   => video_decoder_0_avalon_decoder_source_endofpacket,   --                      .endofpacket
			stream_out_valid         => video_decoder_0_avalon_decoder_source_valid,         --                      .valid
			stream_out_data          => video_decoder_0_avalon_decoder_source_data,          --                      .data
			PIXEL_CLK                => video_in_decoder_PIXEL_CLK,                          --    external_interface.export
			LINE_VALID               => video_in_decoder_LINE_VALID,                         --                      .export
			FRAME_VALID              => video_in_decoder_FRAME_VALID,                        --                      .export
			pixel_clk_reset          => video_in_decoder_pixel_clk_reset,                    --                      .export
			PIXEL_DATA               => video_in_decoder_PIXEL_DATA                          --                      .export
		);

	video_dma_controller : component soc_video_system_video_dma_controller
		port map (
			clk                  => altpll_0_c0_clk,                                                            --                      clk.clk
			reset                => rst_controller_001_reset_out_reset,                                         --                    reset.reset
			stream_data          => video_stream_router_1_avalon_stream_router_source_data,                     --          avalon_dma_sink.data
			stream_startofpacket => video_stream_router_1_avalon_stream_router_source_startofpacket,            --                         .startofpacket
			stream_endofpacket   => video_stream_router_1_avalon_stream_router_source_endofpacket,              --                         .endofpacket
			stream_valid         => video_stream_router_1_avalon_stream_router_source_valid,                    --                         .valid
			stream_ready         => video_stream_router_1_avalon_stream_router_source_ready,                    --                         .ready
			slave_address        => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_address,    -- avalon_dma_control_slave.address
			slave_byteenable     => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_byteenable, --                         .byteenable
			slave_read           => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_read,       --                         .read
			slave_write          => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_write,      --                         .write
			slave_writedata      => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_writedata,  --                         .writedata
			slave_readdata       => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_readdata,   --                         .readdata
			master_address       => video_dma_controller_avalon_dma_master_address,                             --        avalon_dma_master.address
			master_waitrequest   => video_dma_controller_avalon_dma_master_waitrequest,                         --                         .waitrequest
			master_write         => video_dma_controller_avalon_dma_master_write,                               --                         .write
			master_writedata     => video_dma_controller_avalon_dma_master_writedata                            --                         .writedata
		);

	video_dual_clock_buffer : component soc_video_system_video_dual_clock_buffer
		port map (
			clk_stream_in            => altpll_0_c0_clk,                                               --         clock_stream_in.clk
			reset_stream_in          => rst_controller_001_reset_out_reset,                            --         reset_stream_in.reset
			clk_stream_out           => video_pll_vga_clk_clk,                                         --        clock_stream_out.clk
			reset_stream_out         => rst_controller_003_reset_out_reset,                            --        reset_stream_out.reset
			stream_in_ready          => video_pixel_rgb_resampler_1_avalon_rgb_source_ready,           --   avalon_dc_buffer_sink.ready
			stream_in_startofpacket  => video_pixel_rgb_resampler_1_avalon_rgb_source_startofpacket,   --                        .startofpacket
			stream_in_endofpacket    => video_pixel_rgb_resampler_1_avalon_rgb_source_endofpacket,     --                        .endofpacket
			stream_in_valid          => video_pixel_rgb_resampler_1_avalon_rgb_source_valid,           --                        .valid
			stream_in_data           => video_pixel_rgb_resampler_1_avalon_rgb_source_data,            --                        .data
			stream_out_ready         => video_dual_clock_buffer_avalon_dc_buffer_source_ready,         -- avalon_dc_buffer_source.ready
			stream_out_startofpacket => video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket, --                        .startofpacket
			stream_out_endofpacket   => video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket,   --                        .endofpacket
			stream_out_valid         => video_dual_clock_buffer_avalon_dc_buffer_source_valid,         --                        .valid
			stream_out_data          => video_dual_clock_buffer_avalon_dc_buffer_source_data           --                        .data
		);

	video_pixel_buffer_dma : component soc_video_system_video_pixel_buffer_dma
		port map (
			clk                  => altpll_0_c0_clk,                                                          --                     clk.clk
			reset                => rst_controller_001_reset_out_reset,                                       --                   reset.reset
			master_readdatavalid => video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,             -- avalon_pixel_dma_master.readdatavalid
			master_waitrequest   => video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,               --                        .waitrequest
			master_address       => video_pixel_buffer_dma_avalon_pixel_dma_master_address,                   --                        .address
			master_arbiterlock   => video_pixel_buffer_dma_avalon_pixel_dma_master_lock,                      --                        .lock
			master_read          => video_pixel_buffer_dma_avalon_pixel_dma_master_read,                      --                        .read
			master_readdata      => video_pixel_buffer_dma_avalon_pixel_dma_master_readdata,                  --                        .readdata
			slave_address        => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address,    --    avalon_control_slave.address
			slave_byteenable     => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable, --                        .byteenable
			slave_read           => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read,       --                        .read
			slave_write          => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write,      --                        .write
			slave_writedata      => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata,  --                        .writedata
			slave_readdata       => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata,   --                        .readdata
			stream_ready         => video_pixel_buffer_dma_avalon_pixel_source_ready,                         --     avalon_pixel_source.ready
			stream_startofpacket => video_pixel_buffer_dma_avalon_pixel_source_startofpacket,                 --                        .startofpacket
			stream_endofpacket   => video_pixel_buffer_dma_avalon_pixel_source_endofpacket,                   --                        .endofpacket
			stream_valid         => video_pixel_buffer_dma_avalon_pixel_source_valid,                         --                        .valid
			stream_data          => video_pixel_buffer_dma_avalon_pixel_source_data                           --                        .data
		);

	video_pixel_rgb_resampler_1 : component soc_video_system_video_pixel_rgb_resampler_1
		port map (
			clk                      => altpll_0_c0_clk,                                             --               clk.clk
			reset                    => rst_controller_001_reset_out_reset,                          --             reset.reset
			stream_in_startofpacket  => avalon_st_adapter_out_0_startofpacket,                       --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => avalon_st_adapter_out_0_endofpacket,                         --                  .endofpacket
			stream_in_valid          => avalon_st_adapter_out_0_valid,                               --                  .valid
			stream_in_ready          => avalon_st_adapter_out_0_ready,                               --                  .ready
			stream_in_data           => avalon_st_adapter_out_0_data,                                --                  .data
			stream_out_ready         => video_pixel_rgb_resampler_1_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => video_pixel_rgb_resampler_1_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_pixel_rgb_resampler_1_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_pixel_rgb_resampler_1_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => video_pixel_rgb_resampler_1_avalon_rgb_source_data           --                  .data
		);

	video_pll : component soc_video_system_video_pll
		port map (
			ref_clk_clk        => clk_clk,                        --      ref_clk.clk
			ref_reset_reset    => rst_controller_reset_out_reset, --    ref_reset.reset
			video_in_clk_clk   => clk_video_clk,                  -- video_in_clk.clk
			vga_clk_clk        => video_pll_vga_clk_clk,          --      vga_clk.clk
			reset_source_reset => video_pll_reset_source_reset    -- reset_source.reset
		);

	video_rgb_resampler : component soc_video_system_video_rgb_resampler
		port map (
			clk                      => altpll_0_c0_clk,                                     --               clk.clk
			reset                    => rst_controller_001_reset_out_reset,                  --             reset.reset
			stream_in_startofpacket  => video_scaler_avalon_scaler_source_startofpacket,     --   avalon_rgb_sink.startofpacket
			stream_in_endofpacket    => video_scaler_avalon_scaler_source_endofpacket,       --                  .endofpacket
			stream_in_valid          => video_scaler_avalon_scaler_source_valid,             --                  .valid
			stream_in_ready          => video_scaler_avalon_scaler_source_ready,             --                  .ready
			stream_in_data           => video_scaler_avalon_scaler_source_data,              --                  .data
			stream_out_ready         => video_rgb_resampler_avalon_rgb_source_ready,         -- avalon_rgb_source.ready
			stream_out_startofpacket => video_rgb_resampler_avalon_rgb_source_startofpacket, --                  .startofpacket
			stream_out_endofpacket   => video_rgb_resampler_avalon_rgb_source_endofpacket,   --                  .endofpacket
			stream_out_valid         => video_rgb_resampler_avalon_rgb_source_valid,         --                  .valid
			stream_out_data          => video_rgb_resampler_avalon_rgb_source_data           --                  .data
		);

	video_scaler : component soc_video_system_video_scaler
		port map (
			clk                      => altpll_0_c0_clk,                                   --                  clk.clk
			reset                    => rst_controller_001_reset_out_reset,                --                reset.reset
			stream_in_startofpacket  => video_clipper_avalon_clipper_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_clipper_avalon_clipper_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_clipper_avalon_clipper_source_valid,         --                     .valid
			stream_in_ready          => video_clipper_avalon_clipper_source_ready,         --                     .ready
			stream_in_data           => video_clipper_avalon_clipper_source_data,          --                     .data
			stream_out_ready         => video_scaler_avalon_scaler_source_ready,           -- avalon_scaler_source.ready
			stream_out_startofpacket => video_scaler_avalon_scaler_source_startofpacket,   --                     .startofpacket
			stream_out_endofpacket   => video_scaler_avalon_scaler_source_endofpacket,     --                     .endofpacket
			stream_out_valid         => video_scaler_avalon_scaler_source_valid,           --                     .valid
			stream_out_data          => video_scaler_avalon_scaler_source_data             --                     .data
		);

	video_scaler_0 : component soc_video_system_video_scaler_0
		port map (
			clk                      => altpll_0_c0_clk,                                          --                  clk.clk
			reset                    => rst_controller_001_reset_out_reset,                       --                reset.reset
			stream_in_startofpacket  => video_pixel_buffer_dma_avalon_pixel_source_startofpacket, --   avalon_scaler_sink.startofpacket
			stream_in_endofpacket    => video_pixel_buffer_dma_avalon_pixel_source_endofpacket,   --                     .endofpacket
			stream_in_valid          => video_pixel_buffer_dma_avalon_pixel_source_valid,         --                     .valid
			stream_in_ready          => video_pixel_buffer_dma_avalon_pixel_source_ready,         --                     .ready
			stream_in_data           => video_pixel_buffer_dma_avalon_pixel_source_data,          --                     .data
			stream_out_ready         => video_scaler_0_avalon_scaler_source_ready,                -- avalon_scaler_source.ready
			stream_out_startofpacket => video_scaler_0_avalon_scaler_source_startofpacket,        --                     .startofpacket
			stream_out_endofpacket   => video_scaler_0_avalon_scaler_source_endofpacket,          --                     .endofpacket
			stream_out_valid         => video_scaler_0_avalon_scaler_source_valid,                --                     .valid
			stream_out_data          => video_scaler_0_avalon_scaler_source_data,                 --                     .data
			stream_out_channel       => video_scaler_0_avalon_scaler_source_channel               --                     .channel
		);

	video_stream_router_0 : component soc_video_system_video_stream_router_0
		port map (
			clk                        => altpll_0_c0_clk,                                                   --                           clk.clk
			reset                      => rst_controller_001_reset_out_reset,                                --                         reset.reset
			stream_in_data             => video_rgb_resampler_avalon_rgb_source_data,                        --     avalon_stream_router_sink.data
			stream_in_startofpacket    => video_rgb_resampler_avalon_rgb_source_startofpacket,               --                              .startofpacket
			stream_in_endofpacket      => video_rgb_resampler_avalon_rgb_source_endofpacket,                 --                              .endofpacket
			stream_in_valid            => video_rgb_resampler_avalon_rgb_source_valid,                       --                              .valid
			stream_in_ready            => video_rgb_resampler_avalon_rgb_source_ready,                       --                              .ready
			stream_out_ready_0         => video_stream_router_0_avalon_stream_router_source_0_ready,         -- avalon_stream_router_source_0.ready
			stream_out_data_0          => video_stream_router_0_avalon_stream_router_source_0_data,          --                              .data
			stream_out_startofpacket_0 => video_stream_router_0_avalon_stream_router_source_0_startofpacket, --                              .startofpacket
			stream_out_endofpacket_0   => video_stream_router_0_avalon_stream_router_source_0_endofpacket,   --                              .endofpacket
			stream_out_valid_0         => video_stream_router_0_avalon_stream_router_source_0_valid,         --                              .valid
			stream_out_ready_1         => video_stream_router_0_avalon_stream_router_source_1_ready,         -- avalon_stream_router_source_1.ready
			stream_out_data_1          => video_stream_router_0_avalon_stream_router_source_1_data,          --                              .data
			stream_out_startofpacket_1 => video_stream_router_0_avalon_stream_router_source_1_startofpacket, --                              .startofpacket
			stream_out_endofpacket_1   => video_stream_router_0_avalon_stream_router_source_1_endofpacket,   --                              .endofpacket
			stream_out_valid_1         => video_stream_router_0_avalon_stream_router_source_1_valid,         --                              .valid
			stream_select              => video_split_export                                                 --            external_interface.export
		);

	video_stream_router_1 : component soc_video_system_video_stream_router_1
		port map (
			clk                       => altpll_0_c0_clk,                                                   --                         clk.clk
			reset                     => rst_controller_001_reset_out_reset,                                --                       reset.reset
			stream_in_data_0          => video_stream_router_0_avalon_stream_router_source_0_data,          -- avalon_stream_router_sink_0.data
			stream_in_startofpacket_0 => video_stream_router_0_avalon_stream_router_source_0_startofpacket, --                            .startofpacket
			stream_in_endofpacket_0   => video_stream_router_0_avalon_stream_router_source_0_endofpacket,   --                            .endofpacket
			stream_in_valid_0         => video_stream_router_0_avalon_stream_router_source_0_valid,         --                            .valid
			stream_in_ready_0         => video_stream_router_0_avalon_stream_router_source_0_ready,         --                            .ready
			stream_in_data_1          => sobel_edge_detector_0_avalon_streaming_source_data,                -- avalon_stream_router_sink_1.data
			stream_in_startofpacket_1 => sobel_edge_detector_0_avalon_streaming_source_startofpacket,       --                            .startofpacket
			stream_in_endofpacket_1   => sobel_edge_detector_0_avalon_streaming_source_endofpacket,         --                            .endofpacket
			stream_in_valid_1         => sobel_edge_detector_0_avalon_streaming_source_valid,               --                            .valid
			stream_in_ready_1         => sobel_edge_detector_0_avalon_streaming_source_ready,               --                            .ready
			stream_select             => video_merge_export,                                                --          external_interface.export
			stream_out_ready          => video_stream_router_1_avalon_stream_router_source_ready,           -- avalon_stream_router_source.ready
			stream_out_data           => video_stream_router_1_avalon_stream_router_source_data,            --                            .data
			stream_out_startofpacket  => video_stream_router_1_avalon_stream_router_source_startofpacket,   --                            .startofpacket
			stream_out_endofpacket    => video_stream_router_1_avalon_stream_router_source_endofpacket,     --                            .endofpacket
			stream_out_valid          => video_stream_router_1_avalon_stream_router_source_valid            --                            .valid
		);

	video_vga_controller : component soc_video_system_video_vga_controller
		port map (
			clk           => video_pll_vga_clk_clk,                                         --                clk.clk
			reset         => rst_controller_003_reset_out_reset,                            --              reset.reset
			data          => video_dual_clock_buffer_avalon_dc_buffer_source_data,          --    avalon_vga_sink.data
			startofpacket => video_dual_clock_buffer_avalon_dc_buffer_source_startofpacket, --                   .startofpacket
			endofpacket   => video_dual_clock_buffer_avalon_dc_buffer_source_endofpacket,   --                   .endofpacket
			valid         => video_dual_clock_buffer_avalon_dc_buffer_source_valid,         --                   .valid
			ready         => video_dual_clock_buffer_avalon_dc_buffer_source_ready,         --                   .ready
			VGA_CLK       => vga_CLK,                                                       -- external_interface.export
			VGA_HS        => vga_HS,                                                        --                   .export
			VGA_VS        => vga_VS,                                                        --                   .export
			VGA_BLANK     => vga_BLANK,                                                     --                   .export
			VGA_SYNC      => vga_SYNC,                                                      --                   .export
			VGA_R         => vga_R,                                                         --                   .export
			VGA_G         => vga_G,                                                         --                   .export
			VGA_B         => vga_B                                                          --                   .export
		);

	mm_interconnect_0 : component soc_video_system_mm_interconnect_0
		port map (
			altpll_0_c0_clk                                              => altpll_0_c0_clk,                                                               --                                          altpll_0_c0.clk
			clk_0_clk_clk                                                => clk_clk,                                                                       --                                            clk_0_clk.clk
			altpll_0_inclk_interface_reset_reset_bridge_in_reset_reset   => rst_controller_reset_out_reset,                                                -- altpll_0_inclk_interface_reset_reset_bridge_in_reset.reset
			fpga_only_master_clk_reset_reset_bridge_in_reset_reset       => rst_controller_001_reset_out_reset,                                            --     fpga_only_master_clk_reset_reset_bridge_in_reset.reset
			video_dma_controller_reset_reset_bridge_in_reset_reset       => rst_controller_001_reset_out_reset,                                            --     video_dma_controller_reset_reset_bridge_in_reset.reset
			fpga_only_master_master_address                              => fpga_only_master_master_address,                                               --                              fpga_only_master_master.address
			fpga_only_master_master_waitrequest                          => fpga_only_master_master_waitrequest,                                           --                                                     .waitrequest
			fpga_only_master_master_byteenable                           => fpga_only_master_master_byteenable,                                            --                                                     .byteenable
			fpga_only_master_master_read                                 => fpga_only_master_master_read,                                                  --                                                     .read
			fpga_only_master_master_readdata                             => fpga_only_master_master_readdata,                                              --                                                     .readdata
			fpga_only_master_master_readdatavalid                        => fpga_only_master_master_readdatavalid,                                         --                                                     .readdatavalid
			fpga_only_master_master_write                                => fpga_only_master_master_write,                                                 --                                                     .write
			fpga_only_master_master_writedata                            => fpga_only_master_master_writedata,                                             --                                                     .writedata
			video_dma_controller_avalon_dma_master_address               => video_dma_controller_avalon_dma_master_address,                                --               video_dma_controller_avalon_dma_master.address
			video_dma_controller_avalon_dma_master_waitrequest           => video_dma_controller_avalon_dma_master_waitrequest,                            --                                                     .waitrequest
			video_dma_controller_avalon_dma_master_write                 => video_dma_controller_avalon_dma_master_write,                                  --                                                     .write
			video_dma_controller_avalon_dma_master_writedata             => video_dma_controller_avalon_dma_master_writedata,                              --                                                     .writedata
			video_pixel_buffer_dma_avalon_pixel_dma_master_address       => video_pixel_buffer_dma_avalon_pixel_dma_master_address,                        --       video_pixel_buffer_dma_avalon_pixel_dma_master.address
			video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest   => video_pixel_buffer_dma_avalon_pixel_dma_master_waitrequest,                    --                                                     .waitrequest
			video_pixel_buffer_dma_avalon_pixel_dma_master_read          => video_pixel_buffer_dma_avalon_pixel_dma_master_read,                           --                                                     .read
			video_pixel_buffer_dma_avalon_pixel_dma_master_readdata      => video_pixel_buffer_dma_avalon_pixel_dma_master_readdata,                       --                                                     .readdata
			video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid => video_pixel_buffer_dma_avalon_pixel_dma_master_readdatavalid,                  --                                                     .readdatavalid
			video_pixel_buffer_dma_avalon_pixel_dma_master_lock          => video_pixel_buffer_dma_avalon_pixel_dma_master_lock,                           --                                                     .lock
			altpll_0_pll_slave_address                                   => mm_interconnect_0_altpll_0_pll_slave_address,                                  --                                   altpll_0_pll_slave.address
			altpll_0_pll_slave_write                                     => mm_interconnect_0_altpll_0_pll_slave_write,                                    --                                                     .write
			altpll_0_pll_slave_read                                      => mm_interconnect_0_altpll_0_pll_slave_read,                                     --                                                     .read
			altpll_0_pll_slave_readdata                                  => mm_interconnect_0_altpll_0_pll_slave_readdata,                                 --                                                     .readdata
			altpll_0_pll_slave_writedata                                 => mm_interconnect_0_altpll_0_pll_slave_writedata,                                --                                                     .writedata
			audio_and_video_config_0_avalon_av_config_slave_address      => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_address,     --      audio_and_video_config_0_avalon_av_config_slave.address
			audio_and_video_config_0_avalon_av_config_slave_write        => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_write,       --                                                     .write
			audio_and_video_config_0_avalon_av_config_slave_read         => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_read,        --                                                     .read
			audio_and_video_config_0_avalon_av_config_slave_readdata     => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_readdata,    --                                                     .readdata
			audio_and_video_config_0_avalon_av_config_slave_writedata    => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_writedata,   --                                                     .writedata
			audio_and_video_config_0_avalon_av_config_slave_byteenable   => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_byteenable,  --                                                     .byteenable
			audio_and_video_config_0_avalon_av_config_slave_waitrequest  => mm_interconnect_0_audio_and_video_config_0_avalon_av_config_slave_waitrequest, --                                                     .waitrequest
			pixel_buffer_s1_address                                      => mm_interconnect_0_pixel_buffer_s1_address,                                     --                                      pixel_buffer_s1.address
			pixel_buffer_s1_write                                        => mm_interconnect_0_pixel_buffer_s1_write,                                       --                                                     .write
			pixel_buffer_s1_read                                         => mm_interconnect_0_pixel_buffer_s1_read,                                        --                                                     .read
			pixel_buffer_s1_readdata                                     => mm_interconnect_0_pixel_buffer_s1_readdata,                                    --                                                     .readdata
			pixel_buffer_s1_writedata                                    => mm_interconnect_0_pixel_buffer_s1_writedata,                                   --                                                     .writedata
			pixel_buffer_s1_byteenable                                   => mm_interconnect_0_pixel_buffer_s1_byteenable,                                  --                                                     .byteenable
			pixel_buffer_s1_readdatavalid                                => mm_interconnect_0_pixel_buffer_s1_readdatavalid,                               --                                                     .readdatavalid
			pixel_buffer_s1_waitrequest                                  => mm_interconnect_0_pixel_buffer_s1_waitrequest,                                 --                                                     .waitrequest
			pixel_buffer_s1_chipselect                                   => mm_interconnect_0_pixel_buffer_s1_chipselect,                                  --                                                     .chipselect
			pixel_onchip_buffer_s1_address                               => mm_interconnect_0_pixel_onchip_buffer_s1_address,                              --                               pixel_onchip_buffer_s1.address
			pixel_onchip_buffer_s1_write                                 => mm_interconnect_0_pixel_onchip_buffer_s1_write,                                --                                                     .write
			pixel_onchip_buffer_s1_readdata                              => mm_interconnect_0_pixel_onchip_buffer_s1_readdata,                             --                                                     .readdata
			pixel_onchip_buffer_s1_writedata                             => mm_interconnect_0_pixel_onchip_buffer_s1_writedata,                            --                                                     .writedata
			pixel_onchip_buffer_s1_chipselect                            => mm_interconnect_0_pixel_onchip_buffer_s1_chipselect,                           --                                                     .chipselect
			pixel_onchip_buffer_s1_clken                                 => mm_interconnect_0_pixel_onchip_buffer_s1_clken,                                --                                                     .clken
			video_dma_controller_avalon_dma_control_slave_address        => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_address,       --        video_dma_controller_avalon_dma_control_slave.address
			video_dma_controller_avalon_dma_control_slave_write          => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_write,         --                                                     .write
			video_dma_controller_avalon_dma_control_slave_read           => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_read,          --                                                     .read
			video_dma_controller_avalon_dma_control_slave_readdata       => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_readdata,      --                                                     .readdata
			video_dma_controller_avalon_dma_control_slave_writedata      => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_writedata,     --                                                     .writedata
			video_dma_controller_avalon_dma_control_slave_byteenable     => mm_interconnect_0_video_dma_controller_avalon_dma_control_slave_byteenable,    --                                                     .byteenable
			video_pixel_buffer_dma_avalon_control_slave_address          => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_address,         --          video_pixel_buffer_dma_avalon_control_slave.address
			video_pixel_buffer_dma_avalon_control_slave_write            => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_write,           --                                                     .write
			video_pixel_buffer_dma_avalon_control_slave_read             => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_read,            --                                                     .read
			video_pixel_buffer_dma_avalon_control_slave_readdata         => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_readdata,        --                                                     .readdata
			video_pixel_buffer_dma_avalon_control_slave_writedata        => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_writedata,       --                                                     .writedata
			video_pixel_buffer_dma_avalon_control_slave_byteenable       => mm_interconnect_0_video_pixel_buffer_dma_avalon_control_slave_byteenable       --                                                     .byteenable
		);

	avalon_st_adapter : component soc_video_system_avalon_st_adapter
		generic map (
			inBitsPerSymbol => 8,
			inUsePackets    => 1,
			inDataWidth     => 8,
			inChannelWidth  => 2,
			inErrorWidth    => 0,
			inUseEmptyPort  => 0,
			inUseValid      => 1,
			inUseReady      => 1,
			inReadyLatency  => 0,
			outDataWidth    => 8,
			outChannelWidth => 0,
			outErrorWidth   => 0,
			outUseEmptyPort => 0,
			outUseValid     => 1,
			outUseReady     => 1,
			outReadyLatency => 0
		)
		port map (
			in_clk_0_clk        => altpll_0_c0_clk,                                   -- in_clk_0.clk
			in_rst_0_reset      => rst_controller_001_reset_out_reset,                -- in_rst_0.reset
			in_0_data           => video_scaler_0_avalon_scaler_source_data,          --     in_0.data
			in_0_valid          => video_scaler_0_avalon_scaler_source_valid,         --         .valid
			in_0_ready          => video_scaler_0_avalon_scaler_source_ready,         --         .ready
			in_0_startofpacket  => video_scaler_0_avalon_scaler_source_startofpacket, --         .startofpacket
			in_0_endofpacket    => video_scaler_0_avalon_scaler_source_endofpacket,   --         .endofpacket
			in_0_channel        => video_scaler_0_avalon_scaler_source_channel,       --         .channel
			out_0_data          => avalon_st_adapter_out_0_data,                      --    out_0.data
			out_0_valid         => avalon_st_adapter_out_0_valid,                     --         .valid
			out_0_ready         => avalon_st_adapter_out_0_ready,                     --         .ready
			out_0_startofpacket => avalon_st_adapter_out_0_startofpacket,             --         .startofpacket
			out_0_endofpacket   => avalon_st_adapter_out_0_endofpacket                --         .endofpacket
		);

	rst_controller : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => fpga_only_master_master_reset_reset, -- reset_in1.reset
			reset_in2      => video_pll_reset_source_reset,        -- reset_in2.reset
			clk            => clk_clk,                             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,      -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_001 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => fpga_only_master_master_reset_reset, -- reset_in1.reset
			reset_in2      => video_pll_reset_source_reset,        -- reset_in2.reset
			clk            => altpll_0_c0_clk,                     --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_002 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "none",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => fpga_only_master_master_reset_reset, -- reset_in1.reset
			reset_in2      => video_pll_reset_source_reset,        -- reset_in2.reset
			clk            => open,                                --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	rst_controller_003 : component altera_reset_controller
		generic map (
			NUM_RESET_INPUTS          => 3,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,             -- reset_in0.reset
			reset_in1      => fpga_only_master_master_reset_reset, -- reset_in1.reset
			reset_in2      => video_pll_reset_source_reset,        -- reset_in2.reset
			clk            => video_pll_vga_clk_clk,               --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset,  -- reset_out.reset
			reset_req      => open,                                -- (terminated)
			reset_req_in0  => '0',                                 -- (terminated)
			reset_req_in1  => '0',                                 -- (terminated)
			reset_req_in2  => '0',                                 -- (terminated)
			reset_in3      => '0',                                 -- (terminated)
			reset_req_in3  => '0',                                 -- (terminated)
			reset_in4      => '0',                                 -- (terminated)
			reset_req_in4  => '0',                                 -- (terminated)
			reset_in5      => '0',                                 -- (terminated)
			reset_req_in5  => '0',                                 -- (terminated)
			reset_in6      => '0',                                 -- (terminated)
			reset_req_in6  => '0',                                 -- (terminated)
			reset_in7      => '0',                                 -- (terminated)
			reset_req_in7  => '0',                                 -- (terminated)
			reset_in8      => '0',                                 -- (terminated)
			reset_req_in8  => '0',                                 -- (terminated)
			reset_in9      => '0',                                 -- (terminated)
			reset_req_in9  => '0',                                 -- (terminated)
			reset_in10     => '0',                                 -- (terminated)
			reset_req_in10 => '0',                                 -- (terminated)
			reset_in11     => '0',                                 -- (terminated)
			reset_req_in11 => '0',                                 -- (terminated)
			reset_in12     => '0',                                 -- (terminated)
			reset_req_in12 => '0',                                 -- (terminated)
			reset_in13     => '0',                                 -- (terminated)
			reset_req_in13 => '0',                                 -- (terminated)
			reset_in14     => '0',                                 -- (terminated)
			reset_req_in14 => '0',                                 -- (terminated)
			reset_in15     => '0',                                 -- (terminated)
			reset_req_in15 => '0'                                  -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_pixel_buffer_s1_read_ports_inv <= not mm_interconnect_0_pixel_buffer_s1_read;

	mm_interconnect_0_pixel_buffer_s1_byteenable_ports_inv <= not mm_interconnect_0_pixel_buffer_s1_byteenable;

	mm_interconnect_0_pixel_buffer_s1_write_ports_inv <= not mm_interconnect_0_pixel_buffer_s1_write;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of soc_video_system
